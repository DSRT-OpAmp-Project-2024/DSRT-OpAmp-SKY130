magic
tech sky130A
magscale 1 2
timestamp 1718401360
<< pwell >>
rect 878 -2152 8246 -1314
<< metal1 >>
rect 5754 2428 7530 2432
rect 748 2426 7530 2428
rect 560 2226 7530 2426
rect 950 1718 1000 2226
rect 1176 1758 1376 2128
rect 1740 1718 1790 2226
rect 1968 1760 2168 2150
rect 950 110 1066 1718
rect 1478 108 1580 1702
rect 1740 112 1856 1718
rect 2268 112 2380 1710
rect 2520 916 2570 2226
rect 3704 998 3758 2226
rect 3704 960 3860 998
rect 3704 926 3758 960
rect 2520 112 2636 916
rect 3446 912 3560 914
rect 3446 124 3570 912
rect 1540 -40 1580 108
rect 1540 -680 1582 -40
rect 2338 -318 2380 112
rect 3438 62 3570 124
rect 3704 114 3822 926
rect 4634 122 4750 914
rect 4634 118 4638 122
rect 4646 114 4750 122
rect 4892 318 4942 2226
rect 5016 644 6378 734
rect 5016 360 5216 644
rect 5280 318 5320 322
rect 4892 120 5016 318
rect 5206 118 5320 318
rect 2656 38 3570 62
rect 3816 46 4624 64
rect 3520 -178 3570 38
rect 3812 20 4624 46
rect 3812 -178 3966 20
rect 3520 -274 3966 -178
rect 3520 -302 3964 -274
rect 4708 -292 4750 114
rect 5208 106 5320 118
rect 1529 -732 1535 -680
rect 1587 -732 1593 -680
rect 1540 -1210 1582 -732
rect 2338 -1210 2382 -318
rect 1104 -1220 1868 -1210
rect 2296 -1212 3072 -1210
rect 1104 -1262 2000 -1220
rect 1104 -1498 1868 -1262
rect 966 -1544 1040 -1542
rect 1960 -1544 2000 -1262
rect 2296 -1254 3200 -1212
rect 2296 -1498 3072 -1254
rect 3160 -1536 3200 -1254
rect 3520 -1218 3570 -302
rect 4708 -504 4752 -292
rect 4618 -704 4818 -504
rect 4708 -1190 4750 -704
rect 5280 -1002 5320 106
rect 6182 -52 6378 644
rect 6182 -78 6384 -52
rect 6180 -278 6384 -78
rect 6182 -534 6384 -278
rect 6182 -822 6382 -534
rect 5280 -1042 5788 -1002
rect 3520 -1258 4400 -1218
rect 4708 -1236 5598 -1190
rect 4708 -1242 5594 -1236
rect 966 -1944 1088 -1544
rect 1898 -1942 2000 -1544
rect 2166 -1940 2278 -1546
rect 3094 -1938 3200 -1536
rect 4362 -1540 4400 -1258
rect 5006 -1462 5096 -1450
rect 5006 -1528 5012 -1462
rect 5082 -1528 5096 -1462
rect 5006 -1530 5096 -1528
rect 3358 -1938 3472 -1540
rect 966 -1950 1040 -1944
rect 966 -2692 1020 -1950
rect 2166 -2692 2220 -1940
rect 3358 -2692 3400 -1938
rect 4284 -1940 4400 -1540
rect 4346 -1942 4400 -1940
rect 4554 -1946 4670 -1544
rect 5556 -1546 5594 -1242
rect 5482 -1940 5594 -1546
rect 5752 -1844 5788 -1042
rect 5928 -1008 6382 -822
rect 5928 -1720 6036 -1008
rect 6144 -1582 6380 -1540
rect 6144 -1660 6180 -1582
rect 5864 -1810 6066 -1720
rect 5752 -1946 5860 -1844
rect 6070 -1946 6136 -1848
rect 6338 -1846 6380 -1582
rect 7088 -1708 7530 2226
rect 6454 -1758 8052 -1708
rect 6454 -1814 8056 -1758
rect 7088 -1828 7530 -1814
rect 6338 -1920 6448 -1846
rect 6340 -1944 6448 -1920
rect 6138 -1946 6180 -1944
rect 8060 -1946 8176 -1842
rect 4554 -1978 4600 -1946
rect 6070 -1948 6180 -1946
rect 4554 -2018 4694 -1978
rect 4554 -2086 4600 -2018
rect 4554 -2692 4602 -2086
rect 8130 -2692 8176 -1946
rect 766 -2696 8710 -2692
rect 574 -2896 8710 -2696
rect 766 -2898 8710 -2896
<< rmetal1 >>
rect 6144 -1848 6180 -1660
rect 6136 -1944 6180 -1848
rect 6136 -1946 6138 -1944
<< via1 >>
rect 1535 -732 1587 -680
rect 5012 -1528 5082 -1462
<< metal2 >>
rect 1535 -680 1587 -674
rect 1587 -727 5069 -685
rect 1535 -738 1587 -732
rect 5027 -1448 5069 -727
rect 5000 -1462 5096 -1448
rect 5000 -1528 5012 -1462
rect 5082 -1528 5096 -1462
rect 5000 -1542 5096 -1528
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM2
timestamp 1718384992
transform 1 0 1476 0 1 -1740
box -596 -410 596 410
use sky130_fd_pr__pfet_01v8_lvt_ZQZ9VD  XM5
timestamp 1718400045
transform 1 0 4230 0 1 515
box -596 -619 596 619
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM6
timestamp 1718384992
transform 1 0 5068 0 1 -1742
box -596 -410 596 410
use sky130_fd_pr__pfet_01v8_lvt_3VR9VM  XM8
timestamp 1718384992
transform 1 0 5116 0 1 217
box -296 -319 296 319
use sky130_fd_pr__nfet_01v8_lvt_FMMQLY  XM9
timestamp 1718384992
transform 1 0 5956 0 1 -1894
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_lvt_FMHZDY  XM10
timestamp 1718384992
transform 1 0 7252 0 1 -1896
box -996 -260 996 260
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM12
timestamp 1718384992
transform 1 0 3878 0 1 -1736
box -596 -410 596 410
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM18
timestamp 1718384992
transform 1 0 2688 0 1 -1738
box -596 -410 596 410
use sky130_fd_pr__pfet_01v8_lvt_ZQZ9VD  XM54
timestamp 1718400045
transform 1 0 3052 0 1 513
box -596 -619 596 619
use sky130_fd_pr__pfet_01v8_lvt_GWPMZG  XML
timestamp 1718384992
transform 1 0 2076 0 1 915
box -396 -1019 396 1019
use sky130_fd_pr__pfet_01v8_lvt_GWPMZG  XMR
timestamp 1718384992
transform 1 0 1300 0 1 913
box -396 -1019 396 1019
<< labels >>
flabel metal1 560 2226 760 2426 0 FreeSans 256 0 0 0 VCC
port 4 nsew
flabel metal1 574 -2896 774 -2696 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 6180 -278 6380 -78 0 FreeSans 256 0 0 0 ADJ
port 3 nsew
flabel metal1 4618 -704 4818 -504 0 FreeSans 256 0 0 0 DIFFOUT
port 0 nsew
flabel metal1 1968 1950 2168 2150 0 FreeSans 256 0 0 0 MINUS
port 1 nsew
flabel metal1 1176 1928 1376 2128 0 FreeSans 256 0 0 0 PLUS
port 2 nsew
<< end >>
