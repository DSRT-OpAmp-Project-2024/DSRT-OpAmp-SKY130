magic
tech sky130A
magscale 1 2
timestamp 1720781306
<< error_s >>
rect 2893 1226 2928 1260
rect 2894 1207 2928 1226
rect 1015 114 1050 148
rect 2208 131 2242 149
rect 1016 95 1050 114
rect 1035 -600 1050 95
rect 1069 61 1104 95
rect 1069 -600 1103 61
rect 1069 -634 1084 -600
rect 2172 -653 2242 131
rect 2172 -689 2225 -653
rect 2913 -706 2928 1207
rect 2947 1173 2982 1207
rect 2947 -706 2981 1173
rect 7049 214 7084 248
rect 7050 195 7084 214
rect 3633 -28 3667 -10
rect 3633 -64 3703 -28
rect 3650 -98 3721 -64
rect 4771 -98 4806 -64
rect 5964 -81 5998 -63
rect 2947 -740 2962 -706
rect 3650 -759 3720 -98
rect 4772 -117 4806 -98
rect 3650 -795 3703 -759
rect 4791 -812 4806 -117
rect 4825 -151 4860 -117
rect 4825 -812 4859 -151
rect 4825 -846 4840 -812
rect 5928 -865 5998 -81
rect 5928 -901 5981 -865
rect 7069 -918 7084 195
rect 7103 161 7138 195
rect 7103 -918 7137 161
rect 8189 -458 8223 -404
rect 7103 -952 7118 -918
rect 8208 -971 8223 -458
rect 8242 -492 8277 -458
rect 8242 -971 8276 -492
rect 8728 -593 8762 -575
rect 8728 -629 8798 -593
rect 8745 -663 8816 -629
rect 8242 -1005 8257 -971
rect 8745 -1024 8815 -663
rect 8745 -1060 8798 -1024
rect 9286 -1077 9301 -629
rect 9320 -1077 9354 -575
rect 9320 -1111 9335 -1077
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM2 ~/DSRT-OpAmp-SKY130
timestamp 1720781306
transform 1 0 1629 0 1 -279
box -596 -410 596 410
use sky130_fd_pr__pfet_01v8_lvt_ZQZ9VD  XM5 ~/DSRT-OpAmp-SKY130
timestamp 1720781306
transform 1 0 7663 0 1 -388
box -596 -619 596 619
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM6
timestamp 1720781306
transform 1 0 4246 0 1 -438
box -596 -410 596 410
use sky130_fd_pr__pfet_01v8_lvt_3VR9VM  XM8 ~/DSRT-OpAmp-SKY130
timestamp 1720781306
transform 1 0 8502 0 1 -741
box -296 -319 296 319
use sky130_fd_pr__nfet_01v8_lvt_FMMQLY  XM9 ~/DSRT-OpAmp-SKY130
timestamp 1720781306
transform 1 0 9041 0 1 -853
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_lvt_FMHZDY  XM10 ~/DSRT-OpAmp-SKY130
timestamp 1720781306
transform 0 1 9544 -1 0 -170
box -996 -260 996 260
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM12
timestamp 1720781306
transform 1 0 5385 0 1 -491
box -596 -410 596 410
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM18
timestamp 1720781306
transform 1 0 490 0 1 -226
box -596 -410 596 410
use sky130_fd_pr__pfet_01v8_lvt_ZQZ9VD  XM54
timestamp 1720781306
transform 1 0 6524 0 1 -335
box -596 -619 596 619
use sky130_fd_pr__pfet_01v8_lvt_GWPMZG  XML ~/DSRT-OpAmp-SKY130
timestamp 1720781306
transform 1 0 3307 0 1 224
box -396 -1019 396 1019
use sky130_fd_pr__pfet_01v8_lvt_GWPMZG  XMR
timestamp 1720781306
transform 1 0 2568 0 1 277
box -396 -1019 396 1019
<< end >>
